module Switch2Led (Sw,Led);
input [9:0] Sw;
output [9:0] Led;
reg [9:0] Led;
always@(Sw)
begin
	Led[9:0] = Sw[9:0];
end
endmodule