// megafunction wizard: %ALTMULT_ACCUM (MAC)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altmult_accum 

// ============================================================
// File Name: altmult_accum0.v
// Megafunction Name(s):
// 			altmult_accum
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 10.1 Build 153 11/29/2010 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altmult_accum0 (
	aclr0,
	clock0,
	dataa,
	datab,
	overflow,
	result);

	input	  aclr0;
	input	  clock0;
	input	[2:0]  dataa;
	input	[2:0]  datab;
	output	  overflow;
	output	[8:0]  result;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  aclr0;
	tri1	  clock0;
	tri0	[2:0]  dataa;
	tri0	[2:0]  datab;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [8:0] sub_wire1;
	wire  overflow = sub_wire0;
	wire [8:0] result = sub_wire1[8:0];

	altmult_accum	altmult_accum_component (
				.aclr0 (aclr0),
				.clock0 (clock0),
				.datab (datab),
				.dataa (dataa),
				.overflow (sub_wire0),
				.result (sub_wire1),
				.accum_is_saturated (),
				.accum_round (1'b0),
				.accum_saturation (1'b0),
				.accum_sload (1'b0),
				.accum_sload_upper_data (1'b0),
				.aclr1 (1'b0),
				.aclr2 (1'b0),
				.aclr3 (1'b0),
				.addnsub (1'b1),
				.clock1 (1'b1),
				.clock2 (1'b1),
				.clock3 (1'b1),
				.coefsel0 (),
				.coefsel1 (),
				.coefsel2 (),
				.coefsel3 (),
				.datac (),
				.ena0 (1'b1),
				.ena1 (1'b1),
				.ena2 (1'b1),
				.ena3 (1'b1),
				.mult_is_saturated (),
				.mult_round (1'b0),
				.mult_saturation (1'b0),
				.scanina ({3{1'b0}}),
				.scaninb ({3{1'b0}}),
				.scanouta (),
				.scanoutb (),
				.signa (1'b0),
				.signb (1'b0),
				.sourcea (1'b0),
				.sourceb (1'b0));
	defparam
		altmult_accum_component.accum_direction = "ADD",
		altmult_accum_component.addnsub_aclr = "UNUSED",
		altmult_accum_component.addnsub_pipeline_aclr = "UNUSED",
		altmult_accum_component.addnsub_pipeline_reg = "CLOCK0",
		altmult_accum_component.addnsub_reg = "CLOCK0",
		altmult_accum_component.dedicated_multiplier_circuitry = "AUTO",
		altmult_accum_component.input_aclr_a = "UNUSED",
		altmult_accum_component.input_aclr_b = "UNUSED",
		altmult_accum_component.input_reg_a = "CLOCK0",
		altmult_accum_component.input_reg_b = "CLOCK0",
		altmult_accum_component.input_source_a = "DATAA",
		altmult_accum_component.input_source_b = "DATAB",
		altmult_accum_component.intended_device_family = "Cyclone III",
		altmult_accum_component.lpm_type = "altmult_accum",
		altmult_accum_component.multiplier_aclr = "UNUSED",
		altmult_accum_component.multiplier_reg = "CLOCK0",
		altmult_accum_component.output_aclr = "ACLR0",
		altmult_accum_component.output_reg = "CLOCK0",
		altmult_accum_component.port_addnsub = "PORT_UNUSED",
		altmult_accum_component.port_output_is_overflow = "PORT_USED",
		altmult_accum_component.port_signa = "PORT_UNUSED",
		altmult_accum_component.port_signb = "PORT_UNUSED",
		altmult_accum_component.representation_a = "UNSIGNED",
		altmult_accum_component.representation_b = "UNSIGNED",
		altmult_accum_component.sign_aclr_a = "UNUSED",
		altmult_accum_component.sign_aclr_b = "UNUSED",
		altmult_accum_component.sign_pipeline_aclr_a = "UNUSED",
		altmult_accum_component.sign_pipeline_aclr_b = "UNUSED",
		altmult_accum_component.sign_pipeline_reg_a = "CLOCK0",
		altmult_accum_component.sign_pipeline_reg_b = "CLOCK0",
		altmult_accum_component.sign_reg_a = "CLOCK0",
		altmult_accum_component.sign_reg_b = "CLOCK0",
		altmult_accum_component.width_a = 3,
		altmult_accum_component.width_b = 3,
		altmult_accum_component.width_result = 9;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACCUM_SLOAD NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_PIPELINE_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG NUMERIC "1"
// Retrieval info: PRIVATE: ACCUM_SLOAD_REG_INDEX NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_ACLR NUMERIC "3"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_PIPELINE_REG NUMERIC "0"
// Retrieval info: PRIVATE: ACCUM_SLOAD_UPPER_DATA_REG NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
// Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "0"
// Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "0"
// Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: EXTRA_MULTIPLIER_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: HAS_MAC STRING "1"
// Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "0"
// Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "1"
// Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: MULT_LATENCY NUMERIC "0"
// Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "1"
// Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "1"
// Retrieval info: PRIVATE: NUM_MULT STRING "1"
// Retrieval info: PRIVATE: OP1 STRING "Add"
// Retrieval info: PRIVATE: OP3 STRING "Add"
// Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
// Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "0"
// Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW NUMERIC "1"
// Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
// Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
// Retrieval info: PRIVATE: REG_OUT NUMERIC "1"
// Retrieval info: PRIVATE: RNFORMAT STRING "9"
// Retrieval info: PRIVATE: RQFORMAT STRING "Q1.30"
// Retrieval info: PRIVATE: RTS_WIDTH STRING "9"
// Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
// Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
// Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
// Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
// Retrieval info: PRIVATE: SIGNA STRING "UNSIGNED"
// Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNA_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB STRING "UNSIGNED"
// Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
// Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
// Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
// Retrieval info: PRIVATE: SIGNB_REG STRING "1"
// Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIDTHA STRING "3"
// Retrieval info: PRIVATE: WIDTHB STRING "3"
// Retrieval info: PRIVATE: WIDTH_UPPER_DATA NUMERIC "1"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ACCUM_DIRECTION STRING "ADD"
// Retrieval info: CONSTANT: ADDNSUB_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_PIPELINE_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: ADDNSUB_PIPELINE_REG STRING "CLOCK0"
// Retrieval info: CONSTANT: ADDNSUB_REG STRING "CLOCK0"
// Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "AUTO"
// Retrieval info: CONSTANT: INPUT_ACLR_A STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_ACLR_B STRING "UNUSED"
// Retrieval info: CONSTANT: INPUT_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: INPUT_SOURCE_A STRING "DATAA"
// Retrieval info: CONSTANT: INPUT_SOURCE_B STRING "DATAB"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_accum"
// Retrieval info: CONSTANT: MULTIPLIER_ACLR STRING "UNUSED"
// Retrieval info: CONSTANT: MULTIPLIER_REG STRING "CLOCK0"
// Retrieval info: CONSTANT: OUTPUT_ACLR STRING "ACLR0"
// Retrieval info: CONSTANT: OUTPUT_REG STRING "CLOCK0"
// Retrieval info: CONSTANT: PORT_ADDNSUB STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_OUTPUT_IS_OVERFLOW STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: REPRESENTATION_A STRING "UNSIGNED"
// Retrieval info: CONSTANT: REPRESENTATION_B STRING "UNSIGNED"
// Retrieval info: CONSTANT: SIGN_ACLR_A STRING "UNUSED"
// Retrieval info: CONSTANT: SIGN_ACLR_B STRING "UNUSED"
// Retrieval info: CONSTANT: SIGN_PIPELINE_ACLR_A STRING "UNUSED"
// Retrieval info: CONSTANT: SIGN_PIPELINE_ACLR_B STRING "UNUSED"
// Retrieval info: CONSTANT: SIGN_PIPELINE_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGN_PIPELINE_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGN_REG_A STRING "CLOCK0"
// Retrieval info: CONSTANT: SIGN_REG_B STRING "CLOCK0"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "3"
// Retrieval info: CONSTANT: WIDTH_B NUMERIC "3"
// Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "9"
// Retrieval info: USED_PORT: aclr0 0 0 0 0 INPUT GND "aclr0"
// Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
// Retrieval info: USED_PORT: dataa 0 0 3 0 INPUT GND "dataa[2..0]"
// Retrieval info: USED_PORT: datab 0 0 3 0 INPUT GND "datab[2..0]"
// Retrieval info: USED_PORT: overflow 0 0 0 0 OUTPUT NODEFVAL "overflow"
// Retrieval info: USED_PORT: result 0 0 9 0 OUTPUT GND "result[8..0]"
// Retrieval info: CONNECT: @aclr0 0 0 0 0 aclr0 0 0 0 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 3 0 dataa 0 0 3 0
// Retrieval info: CONNECT: @datab 0 0 3 0 datab 0 0 3 0
// Retrieval info: CONNECT: overflow 0 0 0 0 @overflow 0 0 0 0
// Retrieval info: CONNECT: result 0 0 9 0 @result 0 0 9 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altmult_accum0_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
